module TB_four_bit_full_adder (
);

    reg     [3:0]   A_i;
    reg     [3:0]   B_i;
    reg             C_i;
    wire    [3:0]   S_o;
    wire            C_o;

module four_bit_full_adder (
    input   [3:0]   A_i,
    input   [3:0]   B_i,
    input           C_i,
    output  [3:0]   S_o,
    output          C_o
);


endmodule